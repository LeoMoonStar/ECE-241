module ALU(input [7:0] A, B, output [15:0]OUT);

assign OUT = A * B;
	
endmodule 